module raudio

@[typedef]
struct C.rAudioProcessor {
}

type CrAudioProcessor = C.rAudioProcessor
