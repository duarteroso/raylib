module rtextures

type CTexture2D = C.Texture
