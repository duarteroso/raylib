module rtextures

enum BlendMode {
	blend_alpha             = 0
	blend_additive
	blend_multiplied
	blend_add_colors
	blend_subtract_colors
	blend_alpha_premultiply
	blend_custom
	blend_custom_separate
}
