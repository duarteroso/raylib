module raudio

@[typedef]
struct C.rAudioBuffer {
}

type CrAudioBuffer = C.rAudioBuffer
