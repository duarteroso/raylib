module rcore

enum PixelFormat {
	pixelformat_uncompressed_grayscale    = 1
	pixelformat_uncompressed_gray_alpha
	pixelformat_uncompressed_r5g6b5
	pixelformat_uncompressed_r8g8b8
	pixelformat_uncompressed_r5g5b5a1
	pixelformat_uncompressed_r4g4b4a4
	pixelformat_uncompressed_r8g8b8a8
	pixelformat_uncompressed_r32
	pixelformat_uncompressed_r32g32b32
	pixelformat_uncompressed_r32g32b32a32
	pixelformat_uncompressed_r16
	pixelformat_uncompressed_r16g16b16
	pixelformat_uncompressed_r16g16b16a16
	pixelformat_compressed_dxt1_rgb
	pixelformat_compressed_dxt1_rgba
	pixelformat_compressed_dxt3_rgba
	pixelformat_compressed_dxt5_rgba
	pixelformat_compressed_etc1_rgb
	pixelformat_compressed_etc2_rgb
	pixelformat_compressed_etc2_eac_rgba
	pixelformat_compressed_pvrt_rgb
	pixelformat_compressed_pvrt_rgba
	pixelformat_compressed_astc_4x4_rgba
	pixelformat_compressed_astc_8x8_rgba
}
