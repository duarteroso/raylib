module rcore

enum MouseButton {
    mouse_button_left    = 0
    mouse_button_right   = 1
    mouse_button_middle  = 2
    mouse_button_side    = 3
    mouse_button_extra   = 4
    mouse_button_forward = 5
    mouse_button_back    = 6
}