module raylib

$if linux {
}

$if windows {
}
	
$if macos {
	#flag -I/usr/local/inlcude/
	#flag -lraylib
}

#include "raylib.h"