module rcore

enum TraceLogLevel {
	log_all     = 0
	log_trace
	log_debug
	log_info
	log_warning
	log_error
	log_fatal
	log_none
}
