module rcore

enum ShaderUniformDataType {
	shader_uniform_float     = 0
	shader_uniform_vec2
	shader_uniform_vec3
	shader_uniform_vec4
	shader_uniform_int
	shader_uniform_ivec2
	shader_uniform_ivec3
	shader_uniform_ivec4
	shader_uniform_sampler2d
}
