module rtextures

type CTextureCubemap = C.Texture
