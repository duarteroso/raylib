module rtextures

enum TextureWrap {
	texture_wrap_repeat        = 0
	texture_wrap_clamp
	texture_wrap_mirror_repeat
	texture_wrap_mirror_clamp
}
