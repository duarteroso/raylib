module rmath

type CQuaternion = C.Vector4
