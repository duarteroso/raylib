module rmath

@[typedef]
struct C.Vector4 {
pub:
	x f32
	y f32
	z f32
	w f32
}

type CVector4 = C.Vector4
