module rmath

@[typedef]
struct C.Vector2 {
pub:
	x f32
	y f32
}

type CVector2 = C.Vector2
