module rocre

enum CameraProjection {
	camera_perspective  = 0
	camera_orthographic
}
