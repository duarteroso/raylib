module rcore

enum CameraMode {
	camera_custom       = 0
	camera_free
	camera_orbital
	camera_first_person
	camera_third_person
}
