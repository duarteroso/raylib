module rtextures

type CRenderTexture2D = C.RenderTexture
