module rmath

@[typedef]
struct C.Vector3 {
pub:
	x f32
	y f32
	z f32
}

type CVector3 = C.Vector3
