module rtext

enum FontType {
	font_default = 0
	font_bitmap
	font_sdf
}
