module rcore

enum NPatchLayout {
	npatch_nine_patch             = 0
	npatch_three_patch_vertical
	npatch_three_patch_horizontal
}
